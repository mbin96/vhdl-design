library IEEE;
use ieee.std_logic_1164.all;
use ieee.std.logic-unsigned.all;

entity test is
    A
